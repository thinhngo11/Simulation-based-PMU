`include "seq_item.sv"
`include "PMU7seq_item.sv"
`include "PMU10seq_item.sv"
`include "sequence.sv"
`include "seq_full_rw.sv"
`include "seq_7bit.sv"
`include "seq_10bit.sv"
`include "seq_rpt_start.sv"
`include "seq_mismatch.sv"
`include "seq_data_override.sv"
`include "seq_directed.sv"
`include "stuck.sv"

`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "PMU7monitor.sv"
`include "PMU10monitor.sv"
`include "PMU7scoreboard.sv"
`include "PMU10scoreboard.sv"
`include "agent.sv"
`include "PMU7agent.sv"
`include "PMU10agent.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "environment.sv"
`include "test.sv"
